`include "/home/samthekiller/Desktop/Harvard Architecture/My_Code/ALU/Carry Save Array Multiplier/hadd.v"
`include "/home/samthekiller/Desktop/Harvard Architecture/My_Code/ALU/Carry Save Array Multiplier/fadd.v"

module multiplier(x,y,out1);
input [15:0] x;
input [15:0] y;
output [31:0] out1;
    wire a[15:0],b[15:0],c[15:0],d[15:0],e[15:0],f[15:0],g[15:0],h[15:0],i[15:0],j[15:0],k[15:0],l[15:0],m[15:0],n[15:0],o[15:0],p[15:0];
    wire carry1[14:0],carry2[14:0],carry3[14:0],carry4[14:0],carry5[14:0],carry6[14:0],carry7[14:0];
    wire carry8[14:0],carry9[14:0],carry10[14:0],carry11[14:0],carry12[14:0],carry13[14:0],carry14[14:0],carry15[14:0],carry16[14:0];
    wire sum1[14:0],sum2[14:0],sum3[14:0],sum4[14:0],sum5[14:0],sum6[14:0],sum7[14:0],sum8[14:0];
    wire sum9[14:0],sum10[14:0],sum11[14:0],sum12[14:0],sum13[14:0],sum14[14:0],sum15[14:0];

    assign a[0]=x[0] & y[0];
    assign a[1]=x[1] & y[0];
    assign a[2]=x[2] & y[0];
    assign a[3]=x[3] & y[0];
    assign a[4]=x[4] & y[0];
    assign a[5]=x[5] & y[0];
    assign a[6]=x[6] & y[0];
    assign a[7]=x[7] & y[0];
    assign a[8]=x[8] & y[0];
    assign a[9]=x[9] & y[0];
    assign a[10]=x[10] & y[0];
    assign a[11]=x[11] & y[0];
    assign a[12]=x[12] & y[0];
    assign a[13]=x[13] & y[0];
    assign a[14]=x[14] & y[0];
    assign a[15]=x[15] & y[0];

    assign b[0]=x[0] & y[1];
    assign b[1]=x[1] & y[1];
    assign b[2]=x[2] & y[1];
    assign b[3]=x[3] & y[1];
    assign b[4]=x[4] & y[1];
    assign b[5]=x[5] & y[1];
    assign b[6]=x[6] & y[1];
    assign b[7]=x[7] & y[1];
    assign b[8]=x[8] & y[1];
    assign b[9]=x[9] & y[1];
    assign b[10]=x[10] & y[1];
    assign b[11]=x[11] & y[1];
    assign b[12]=x[12] & y[1];
    assign b[13]=x[13] & y[1];
    assign b[14]=x[14] & y[1];
    assign b[15]=x[15] & y[1];

    assign c[0]=x[0] & y[2];
    assign c[1]=x[1] & y[2];
    assign c[2]=x[2] & y[2];
    assign c[3]=x[3] & y[2];
    assign c[4]=x[4] & y[2];
    assign c[5]=x[5] & y[2];
    assign c[6]=x[6] & y[2];
    assign c[7]=x[7] & y[2];
    assign c[8]=x[8] & y[2];
    assign c[9]=x[9] & y[2];
    assign c[10]=x[10] & y[2];
    assign c[11]=x[11] & y[2];
    assign c[12]=x[12] & y[2];
    assign c[13]=x[13] & y[2];
    assign c[14]=x[14] & y[2];
    assign c[15]=x[15] & y[2];

    assign d[0]=x[0] & y[3];
    assign d[1]=x[1] & y[3];
    assign d[2]=x[2] & y[3];
    assign d[3]=x[3] & y[3];
    assign d[4]=x[4] & y[3];
    assign d[5]=x[5] & y[3];
    assign d[6]=x[6] & y[3];
    assign d[7]=x[7] & y[3];
    assign d[8]=x[8] & y[3];
    assign d[9]=x[9] & y[3];
    assign d[10]=x[10] & y[3];
    assign d[11]=x[11] & y[3];
    assign d[12]=x[12] & y[3];
    assign d[13]=x[13] & y[3];
    assign d[14]=x[14] & y[3];
    assign d[15]=x[15] & y[3];

    assign e[0]=x[0] & y[4];
    assign e[1]=x[1] & y[4];
    assign e[2]=x[2] & y[4];
    assign e[3]=x[3] & y[4];
    assign e[4]=x[4] & y[4];
    assign e[5]=x[5] & y[4];
    assign e[6]=x[6] & y[4];
    assign e[7]=x[7] & y[4];
    assign e[8]=x[8] & y[4];
    assign e[9]=x[9] & y[4];
    assign e[10]=x[10] & y[4];
    assign e[11]=x[11] & y[4];
    assign e[12]=x[12] & y[4];
    assign e[13]=x[13] & y[4];
    assign e[14]=x[14] & y[4];
    assign e[15]=x[15] & y[4];

    assign f[0]=x[0] & y[5];
    assign f[1]=x[1] & y[5];
    assign f[2]=x[2] & y[5];
    assign f[3]=x[3] & y[5];
    assign f[4]=x[4] & y[5];
    assign f[5]=x[5] & y[5];
    assign f[6]=x[6] & y[5];
    assign f[7]=x[7] & y[5];
    assign f[8]=x[8] & y[5];
    assign f[9]=x[9] & y[5];
    assign f[10]=x[10] & y[5];
    assign f[11]=x[11] & y[5];
    assign f[12]=x[12] & y[5];
    assign f[13]=x[13] & y[5];
    assign f[14]=x[14] & y[5];
    assign f[15]=x[15] & y[5];

    assign g[0]=x[0] & y[6];
    assign g[1]=x[1] & y[6];
    assign g[2]=x[2] & y[6];
    assign g[3]=x[3] & y[6];
    assign g[4]=x[4] & y[6];
    assign g[5]=x[5] & y[6];
    assign g[6]=x[6] & y[6];
    assign g[7]=x[7] & y[6];
    assign g[8]=x[8] & y[6];
    assign g[9]=x[9] & y[6];
    assign g[10]=x[10] & y[6];
    assign g[11]=x[11] & y[6];
    assign g[12]=x[12] & y[6];
    assign g[13]=x[13] & y[6];
    assign g[14]=x[14] & y[6];
    assign g[15]=x[15] & y[6];

    assign h[0]=x[0] & y[7];
    assign h[1]=x[1] & y[7];
    assign h[2]=x[2] & y[7];
    assign h[3]=x[3] & y[7];
    assign h[4]=x[4] & y[7];
    assign h[5]=x[5] & y[7];
    assign h[6]=x[6] & y[7];
    assign h[7]=x[7] & y[7];
    assign h[8]=x[8] & y[7];
    assign h[9]=x[9] & y[7];
    assign h[10]=x[10] & y[7];
    assign h[11]=x[11] & y[7];
    assign h[12]=x[12] & y[7];
    assign h[13]=x[13] & y[7];
    assign h[14]=x[14] & y[7];
    assign h[15]=x[15] & y[7];

    assign i[0]=x[0] & y[8];
    assign i[1]=x[1] & y[8];
    assign i[2]=x[2] & y[8];
    assign i[3]=x[3] & y[8];
    assign i[4]=x[4] & y[8];
    assign i[5]=x[5] & y[8];
    assign i[6]=x[6] & y[8];
    assign i[7]=x[7] & y[8];
    assign i[8]=x[8] & y[8];
    assign i[9]=x[9] & y[8];
    assign i[10]=x[10] & y[8];
    assign i[11]=x[11] & y[8];
    assign i[12]=x[12] & y[8];
    assign i[13]=x[12] & y[8];
    assign i[14]=x[12] & y[8];
    assign i[15]=x[12] & y[8];

    assign j[0]=x[0] & y[9];
    assign j[1]=x[1] & y[9];
    assign j[2]=x[2] & y[9];
    assign j[3]=x[3] & y[9];
    assign j[4]=x[4] & y[9];
    assign j[5]=x[5] & y[9];
    assign j[6]=x[6] & y[9];
    assign j[7]=x[7] & y[9];
    assign j[8]=x[8] & y[9];
    assign j[9]=x[9] & y[9];
    assign j[10]=x[10] & y[9];
    assign j[11]=x[11] & y[9];
    assign j[12]=x[12] & y[9];
    assign j[13]=x[13] & y[9];
    assign j[14]=x[14] & y[9];
    assign j[15]=x[15] & y[9];

    assign k[0]=x[0] & y[10];
    assign k[1]=x[1] & y[10];
    assign k[2]=x[2] & y[10];
    assign k[3]=x[3] & y[10];
    assign k[4]=x[4] & y[10];
    assign k[5]=x[5] & y[10];
    assign k[6]=x[6] & y[10];
    assign k[7]=x[7] & y[10];
    assign k[8]=x[8] & y[10];
    assign k[9]=x[9] & y[10];
    assign k[10]=x[10] & y[10];
    assign k[11]=x[11] & y[10];
    assign k[12]=x[12] & y[10];
    assign k[13]=x[13] & y[10];
    assign k[14]=x[14] & y[10];
    assign k[15]=x[15] & y[10];

    assign l[0]=x[0] & y[11];
    assign l[1]=x[1] & y[11];
    assign l[2]=x[2] & y[11];
    assign l[3]=x[3] & y[11];
    assign l[4]=x[4] & y[11];
    assign l[5]=x[5] & y[11];
    assign l[6]=x[6] & y[11];
    assign l[7]=x[7] & y[11];
    assign l[8]=x[8] & y[11];
    assign l[9]=x[9] & y[11];
    assign l[10]=x[10] & y[11];
    assign l[11]=x[11] & y[11];
    assign l[12]=x[12] & y[11];
    assign l[13]=x[13] & y[11];
    assign l[14]=x[14] & y[11];
    assign l[15]=x[15] & y[11];

    assign m[0]=x[0] & y[12];
    assign m[1]=x[1] & y[12];
    assign m[2]=x[2] & y[12];
    assign m[3]=x[3] & y[12];
    assign m[4]=x[4] & y[12];
    assign m[5]=x[5] & y[12];
    assign m[6]=x[6] & y[12];
    assign m[7]=x[7] & y[12];
    assign m[8]=x[8] & y[12];
    assign m[9]=x[9] & y[12];
    assign m[10]=x[10] & y[12];
    assign m[11]=x[11] & y[12];
    assign m[12]=x[12] & y[12];
    assign m[13]=x[13] & y[12];
    assign m[14]=x[14] & y[12];
    assign m[15]=x[15] & y[12];

    assign n[0]=x[0] & y[13];
    assign n[1]=x[1] & y[13];
    assign n[2]=x[2] & y[13];
    assign n[3]=x[3] & y[13];
    assign n[4]=x[4] & y[13];
    assign n[5]=x[5] & y[13];
    assign n[6]=x[6] & y[13];
    assign n[7]=x[7] & y[13];
    assign n[8]=x[8] & y[13];
    assign n[9]=x[9] & y[13];
    assign n[10]=x[10] & y[13];
    assign n[11]=x[11] & y[13];
    assign n[12]=x[12] & y[13];
    assign n[13]=x[13] & y[13];
    assign n[14]=x[14] & y[13];
    assign n[15]=x[15] & y[13];

    assign o[0]=x[0] & y[14];
    assign o[1]=x[1] & y[14];
    assign o[2]=x[2] & y[14];
    assign o[3]=x[3] & y[14];
    assign o[4]=x[4] & y[14];
    assign o[5]=x[5] & y[14];
    assign o[6]=x[6] & y[14];
    assign o[7]=x[7] & y[14];
    assign o[8]=x[8] & y[14];
    assign o[9]=x[9] & y[14];
    assign o[10]=x[10] & y[14];
    assign o[11]=x[11] & y[14];
    assign o[12]=x[12] & y[14];
    assign o[13]=x[13] & y[14];
    assign o[14]=x[14] & y[14];
    assign o[15]=x[15] & y[14];

    assign p[0]=x[0] & y[15];
    assign p[1]=x[1] & y[15];
    assign p[2]=x[2] & y[15];
    assign p[3]=x[3] & y[15];
    assign p[4]=x[4] & y[15];
    assign p[5]=x[5] & y[15];
    assign p[6]=x[6] & y[15];
    assign p[7]=x[7] & y[15];
    assign p[8]=x[8] & y[15];
    assign p[9]=x[9] & y[15];
    assign p[10]=x[10] & y[15];
    assign p[11]=x[11] & y[15];
    assign p[12]=x[12] & y[15];
    assign p[13]=x[13] & y[15];
    assign p[14]=x[14] & y[15];
    assign p[15]=x[15] & y[15];



    assign out1[0]=a[0];

    half_adder h11(a[1],b[0],out1[1],carry1[0]);

    full_adder f11(a[2],b[1],c[0],sum1[0],carry1[1]);
    half_adder h1_1(sum1[0],carry1[0],out1[2],carry2[0]);

    full_adder f21(a[3],b[2],c[1],sum1[1],carry1[2]);
    full_adder f22(d[0],sum1[1],carry1[1],sum2[0],carry2[1]);
    half_adder h2_2(sum2[0],carry2[0],out1[3],carry3[0]);

    full_adder f31(a[4],b[3],c[2],sum1[2],carry1[3]);
    full_adder f32(d[1],sum1[2],carry1[2],sum2[1],carry2[2]);
    full_adder f33(e[0],sum2[1],carry2[1],sum3[0],carry3[1]);
    half_adder h3_3(sum3[0],carry3[0],out1[4],carry4[0]);

    full_adder f41(a[5],b[4],c[3],sum1[3],carry1[4]);
    full_adder f42(d[2],sum1[3],carry1[3],sum2[2],carry2[3]);
    full_adder f43(e[1],sum2[2],carry2[2],sum3[1],carry3[2]);
    full_adder f44(f[0],sum3[1],carry3[1],sum4[0],carry4[1]);
    half_adder h4_4(sum4[0],carry4[0],out1[5],carry5[0]);

    full_adder f51(a[6],b[5],c[4],sum1[4],carry1[5]);
    full_adder f52(d[3],sum1[4],carry1[4],sum2[3],carry2[4]);
    full_adder f53(e[2],sum2[3],carry2[3],sum3[2],carry3[3]);
    full_adder f54(f[1],sum3[2],carry3[2],sum4[1],carry4[2]);
    full_adder f55(g[0],sum4[1],carry4[1],sum5[0],carry5[1]);
    half_adder h5_5(sum5[0],carry5[0],out1[6],carry6[0]);

    full_adder f61(a[7],b[6],c[5],sum1[5],carry1[6]);
    full_adder f62(d[4],sum1[5],carry1[5],sum2[4],carry2[5]);
    full_adder f63(e[3],sum2[4],carry2[4],sum3[3],carry3[4]);
    full_adder f64(f[2],sum3[3],carry3[3],sum4[2],carry4[3]);
    full_adder f65(g[1],sum4[2],carry4[2],sum5[1],carry5[2]);
    full_adder f66(h[0],sum5[1],carry5[1],sum6[0],carry6[1]);
    half_adder h6_6(sum6[0],carry6[0],out1[7],carry7[0]);

    full_adder f71(a[8],b[7],c[6],sum1[6],carry1[7]);
    full_adder f72(d[5],sum1[6],carry1[6],sum2[5],carry2[6]);
    full_adder f73(e[4],sum2[5],carry2[5],sum3[4],carry3[5]);
    full_adder f74(f[3],sum3[4],carry3[4],sum4[3],carry4[4]);
    full_adder f75(g[2],sum4[3],carry4[3],sum5[2],carry5[3]);
    full_adder f76(h[1],sum5[2],carry5[2],sum6[1],carry6[2]);
    full_adder f77(i[0],sum6[1],carry6[1],sum7[0],carry7[1]);
    half_adder h7_7(sum7[0],carry7[0],out1[8],carry8[0]);

    full_adder f81(a[9],b[8],c[7],sum1[7],carry1[8]);
    full_adder f82(d[6],sum1[7],carry1[7],sum2[6],carry2[7]);
    full_adder f83(e[5],sum2[6],carry2[6],sum3[5],carry3[6]);
    full_adder f84(f[4],sum3[5],carry3[5],sum4[4],carry4[5]);
    full_adder f85(g[3],sum4[4],carry4[4],sum5[3],carry5[4]);
    full_adder f86(h[2],sum5[3],carry5[3],sum6[2],carry6[3]);
    full_adder f87(i[1],sum6[2],carry6[2],sum7[1],carry7[2]);
    full_adder f88(j[0],sum7[1],carry7[1],sum8[0],carry8[1]);
    half_adder h8_8(sum8[0],carry8[0],out1[9],carry9[0]);

    full_adder f91(a[10],b[9],c[8],sum1[8],carry1[9]);
    full_adder f92(d[7],sum1[8],carry1[8],sum2[7],carry2[8]);
    full_adder f93(e[6],sum2[7],carry2[7],sum3[6],carry3[7]);
    full_adder f94(f[5],sum3[6],carry3[6],sum4[5],carry4[6]);
    full_adder f95(g[4],sum4[5],carry4[5],sum5[4],carry5[5]);
    full_adder f96(h[3],sum5[4],carry5[4],sum6[3],carry6[4]);
    full_adder f97(i[2],sum6[3],carry6[3],sum7[2],carry7[3]);
    full_adder f98(j[1],sum7[2],carry7[2],sum8[1],carry8[2]);
    full_adder f99(k[0],sum8[1],carry8[1],sum9[0],carry9[1]);
    half_adder h9_9(sum9[0],carry9[0],out1[10],carry10[0]);

    full_adder f10_1(a[11],b[10],c[9],sum1[9],carry1[10]);
    full_adder f10_2(d[8],sum1[9],carry1[9],sum2[8],carry2[9]);
    full_adder f10_3(e[7],sum2[8],carry2[8],sum3[7],carry3[8]);
    full_adder f10_4(f[6],sum3[7],carry3[7],sum4[6],carry4[7]);
    full_adder f10_5(g[5],sum4[6],carry4[6],sum5[5],carry5[6]);
    full_adder f10_6(h[4],sum5[5],carry5[5],sum6[4],carry6[5]);
    full_adder f10_7(i[3],sum6[4],carry6[4],sum7[3],carry7[4]);
    full_adder f10_8(j[2],sum7[3],carry7[3],sum8[2],carry8[3]);
    full_adder f10_9(k[1],sum8[2],carry8[2],sum9[1],carry9[2]);
    full_adder f10_10(l[0],sum9[1],carry9[1],sum10[0],carry10[1]);
    half_adder h10_10(sum10[0],carry10[0],out1[11],carry11[0]);

    full_adder f11_1(a[12],b[11],c[10],sum1[10],carry1[11]);
    full_adder f11_2(d[9],sum1[10],carry1[10],sum2[9],carry2[10]);
    full_adder f11_3(e[8],sum2[9],carry2[9],sum3[8],carry3[9]);
    full_adder f11_4(f[7],sum3[8],carry3[8],sum4[7],carry4[8]);
    full_adder f11_5(g[6],sum4[7],carry4[7],sum5[6],carry5[7]);
    full_adder f11_6(h[5],sum5[6],carry5[6],sum6[5],carry6[6]);
    full_adder f11_7(i[4],sum6[5],carry6[5],sum7[4],carry7[5]);
    full_adder f11_8(j[3],sum7[4],carry7[4],sum8[3],carry8[4]);
    full_adder f11_9(k[2],sum8[3],carry8[3],sum9[2],carry9[3]);
    full_adder f11_10(l[1],sum9[2],carry9[2],sum10[1],carry10[2]);
    full_adder f11_11(m[0],sum10[1],carry10[1],sum11[0],carry11[1]);
    half_adder h11_11(sum11[0],carry11[0],out1[12],carry12[0]);

    full_adder f12_1(a[13],b[12],c[11],sum1[11],carry1[12]);
    full_adder f12_2(d[10],sum1[11],carry1[11],sum2[10],carry2[11]);
    full_adder f12_3(e[9],sum2[10],carry2[10],sum3[9],carry3[10]);
    full_adder f12_4(f[8],sum3[9],carry3[9],sum4[8],carry4[9]);
    full_adder f12_5(g[7],sum4[8],carry4[8],sum5[7],carry5[8]);
    full_adder f12_6(h[6],sum5[7],carry5[7],sum6[6],carry6[7]);
    full_adder f12_7(i[5],sum6[6],carry6[6],sum7[5],carry7[6]);
    full_adder f12_8(j[4],sum7[5],carry7[5],sum8[4],carry8[5]);
    full_adder f12_9(k[3],sum8[4],carry8[4],sum9[3],carry9[4]);
    full_adder f12_10(l[2],sum9[3],carry9[3],sum10[2],carry10[3]);
    full_adder f12_11(m[1],sum10[2],carry10[2],sum11[1],carry11[2]);
    full_adder f12_12(n[0],sum11[1],carry11[1],sum12[0],carry12[1]);
    half_adder h12_12(sum12[0],carry12[0],out1[13],carry13[0]);

    full_adder f13_1(a[14],b[13],c[12],sum1[12],carry1[13]);
    full_adder f13_2(d[11],sum1[12],carry1[12],sum2[11],carry2[12]);
    full_adder f13_3(e[10],sum2[11],carry2[11],sum3[10],carry3[11]);
    full_adder f13_4(f[9],sum3[10],carry3[10],sum4[9],carry4[10]);
    full_adder f13_5(g[8],sum4[9],carry4[9],sum5[8],carry5[9]);
    full_adder f13_6(h[7],sum5[8],carry5[8],sum6[7],carry6[8]);
    full_adder f13_7(i[6],sum6[7],carry6[7],sum7[6],carry7[7]);
    full_adder f13_8(j[5],sum7[6],carry7[6],sum8[5],carry8[6]);
    full_adder f13_9(k[4],sum8[5],carry8[5],sum9[4],carry9[5]);
    full_adder f13_10(l[3],sum9[4],carry9[4],sum10[3],carry10[4]);
    full_adder f13_11(m[2],sum10[3],carry10[3],sum11[2],carry11[3]);
    full_adder f13_12(n[1],sum11[2],carry11[2],sum12[1],carry12[2]);
    full_adder f13_13(o[0],sum12[1],carry12[1],sum13[0],carry13[1]);
    half_adder h13_13(sum13[0],carry13[0],out1[14],carry14[0]);

    full_adder f14_1(a[15],b[14],c[13],sum1[13],carry1[14]);
    full_adder f14_2(d[12],sum1[13],carry1[13],sum2[12],carry2[13]);
    full_adder f14_3(e[11],sum2[12],carry2[12],sum3[11],carry3[12]);
    full_adder f14_4(f[10],sum3[11],carry3[11],sum4[10],carry4[11]);
    full_adder f14_5(g[9],sum4[10],carry4[10],sum5[9],carry5[10]);
    full_adder f14_6(h[8],sum5[9],carry5[9],sum6[8],carry6[9]);
    full_adder f14_7(i[7],sum6[8],carry6[8],sum7[7],carry7[8]);
    full_adder f14_8(j[6],sum7[7],carry7[7],sum8[6],carry8[7]);
    full_adder f14_9(k[5],sum8[6],carry8[6],sum9[5],carry9[6]);
    full_adder f14_10(l[4],sum9[5],carry9[5],sum10[4],carry10[5]);
    full_adder f14_11(m[3],sum10[4],carry10[4],sum11[3],carry11[4]);
    full_adder f14_12(n[2],sum11[3],carry11[3],sum12[2],carry12[3]);
    full_adder f14_13(o[1],sum12[2],carry12[2],sum13[1],carry13[2]);
    full_adder f14_14(p[0],sum13[1],carry13[1],sum14[0],carry14[1]);
    half_adder h14_14(sum14[0],carry14[0],out1[15],carry15[0]);





    full_adder f14_1_(b[15],c[14],carry1[14],sum2[13],carry2[14]);
    full_adder f14_2_(d[13],sum2[13],carry2[13],sum3[12],carry3[13]);
    full_adder f14_3_(e[12],sum3[12],carry3[12],sum4[11],carry4[12]);
    full_adder f14_4_(f[11],sum4[11],carry4[11],sum5[10],carry5[11]);
    full_adder f14_5_(g[10],sum5[10],carry5[10],sum6[9],carry6[10]);
    full_adder f14_6_(h[9],sum6[9],carry6[9],sum7[8],carry7[9]);
    full_adder f14_7_(i[8],sum7[8],carry7[8],sum8[7],carry8[8]);
    full_adder f14_8_(j[7],sum8[7],carry8[7],sum9[6],carry9[7]);
    full_adder f14_9_(k[6],sum9[6],carry9[6],sum10[5],carry10[6]);
    full_adder f14_10_(l[5],sum10[5],carry10[5],sum11[4],carry11[5]);
    full_adder f14_11_(m[4],sum11[4],carry11[4],sum12[3],carry12[4]);
    full_adder f14_12_(n[3],sum12[3],carry12[3],sum13[2],carry13[3]);
    full_adder f14_13_(o[2],sum13[2],carry13[2],sum14[1],carry14[2]);
    full_adder f14_14_(p[1],sum14[1],carry14[1],sum15[0],carry15[1]);
    half_adder h14_14_(sum15[0],carry15[0],out1[16],carry16[0]);

    full_adder f113_1(c[15],d[14],carry2[14],sum3[13],carry3[14]);
    full_adder f113_2(e[13],sum3[13],carry3[13],sum4[12],carry4[13]);
    full_adder f113_3(f[12],sum4[12],carry4[12],sum5[11],carry5[12]);
    full_adder f113_4(g[11],sum5[11],carry5[11],sum6[10],carry6[11]);
    full_adder f113_5(h[10],sum6[10],carry6[10],sum7[9],carry7[10]);
    full_adder f113_6(i[9],sum7[9],carry7[9],sum8[8],carry8[9]);
    full_adder f113_7(j[8],sum8[8],carry8[8],sum9[7],carry9[8]);
    full_adder f113_8(k[7],sum9[7],carry9[7],sum10[6],carry10[7]);
    full_adder f113_9(l[6],sum10[6],carry10[6],sum11[5],carry11[6]);
    full_adder f113_10(m[5],sum11[5],carry11[5],sum12[4],carry12[5]);
    full_adder f113_11(n[4],sum12[4],carry12[4],sum13[3],carry13[4]);
    full_adder f113_12(o[3],sum13[3],carry13[3],sum14[2],carry14[3]);
    full_adder f113_13(p[2],sum14[2],carry14[2],sum15[1],carry15[2]);
    full_adder f113_14(sum15[1],carry15[1],carry16[0],out1[17],carry16[1]);

    full_adder f112_1(d[15],e[14],carry3[14],sum4[13],carry4[14]);
    full_adder f112_2(f[13],sum4[13],carry4[13],sum5[12],carry5[13]);
    full_adder f112_3(g[12],sum5[12],carry5[12],sum6[11],carry6[12]);
    full_adder f112_4(h[11],sum6[11],carry6[11],sum7[10],carry7[11]);
    full_adder f112_5(i[10],sum7[10],carry7[10],sum8[9],carry8[10]);
    full_adder f112_6(j[9],sum8[9],carry8[9],sum9[8],carry9[9]);
    full_adder f112_7(k[8],sum9[8],carry9[8],sum10[7],carry10[8]);
    full_adder f112_8(l[7],sum10[7],carry10[7],sum11[6],carry11[7]);
    full_adder f112_9(m[6],sum11[6],carry11[6],sum12[5],carry12[6]);
    full_adder f112_10(n[5],sum12[5],carry12[5],sum13[4],carry13[5]);
    full_adder f112_11(o[4],sum13[4],carry13[4],sum14[3],carry14[4]);
    full_adder f112_12(p[3],sum14[3],carry14[3],sum15[2],carry15[3]);
    full_adder f112_13(sum15[2],carry15[2],carry16[1],out1[18],carry16[2]);

    full_adder f111_1(e[15],f[14],carry4[14],sum5[13],carry5[14]);
    full_adder f111_2(g[13],sum5[13],carry5[13],sum6[12],carry6[13]);
    full_adder f111_3(h[12],sum6[12],carry6[12],sum7[11],carry7[12]);
    full_adder f111_4(i[11],sum7[11],carry7[11],sum8[10],carry8[11]);
    full_adder f111_5(j[10],sum8[10],carry8[10],sum9[9],carry9[10]);
    full_adder f111_6(k[9],sum9[9],carry9[9],sum10[8],carry10[9]);
    full_adder f111_7(l[8],sum10[8],carry10[8],sum11[7],carry11[8]);
    full_adder f111_8(m[7],sum11[7],carry11[7],sum12[6],carry12[7]);
    full_adder f111_9(n[6],sum12[6],carry12[6],sum13[5],carry13[6]);
    full_adder f111_10(o[5],sum13[5],carry13[5],sum14[4],carry14[5]);
    full_adder f111_11(p[4],sum14[4],carry14[4],sum15[3],carry15[4]);
    full_adder f111_12(sum15[3],carry15[3],carry16[2],out1[19],carry16[3]);

    full_adder f110_1(f[15],g[14],carry5[14],sum6[13],carry6[14]);
    full_adder f110_2(h[13],sum6[13],carry6[13],sum7[12],carry7[13]);
    full_adder f110_3(i[12],sum7[12],carry7[12],sum8[11],carry8[12]);
    full_adder f110_4(j[11],sum8[11],carry8[11],sum9[10],carry9[11]);
    full_adder f110_5(k[10],sum9[10],carry9[10],sum10[9],carry10[10]);
    full_adder f110_6(l[9],sum10[9],carry10[9],sum11[8],carry11[9]);
    full_adder f110_7(m[8],sum11[8],carry11[8],sum12[7],carry12[8]);
    full_adder f110_8(n[7],sum12[7],carry12[7],sum13[6],carry13[7]);
    full_adder f110_9(o[6],sum13[6],carry13[6],sum14[5],carry14[6]);
    full_adder f110_10(p[5],sum14[5],carry14[5],sum15[4],carry15[5]);
    full_adder f110_11(sum15[4],carry15[4],carry16[3],out1[20],carry16[4]);

    full_adder f9_1(g[15],h[14],carry6[14],sum7[13],carry7[14]);
    full_adder f9_2(i[13],sum7[13],carry7[13],sum8[12],carry8[13]);
    full_adder f9_3(j[12],sum8[12],carry8[12],sum9[11],carry9[12]);
    full_adder f9_4(k[11],sum9[11],carry9[11],sum10[10],carry10[11]);
    full_adder f9_5(l[10],sum10[10],carry10[10],sum11[9],carry11[10]);
    full_adder f9_6(m[9],sum11[9],carry11[9],sum12[8],carry12[9]);
    full_adder f9_7(n[8],sum12[8],carry12[8],sum13[7],carry13[8]);
    full_adder f9_8(o[7],sum13[7],carry13[7],sum14[6],carry14[7]);
    full_adder f9_9(p[6],sum14[6],carry14[6],sum15[5],carry15[6]);
    full_adder f9_10(sum15[5],carry15[5],carry16[4],out1[21],carry16[5]);

    full_adder f8_1(h[15],i[14],carry7[14],sum8[13],carry8[14]);
    full_adder f8_2(j[13],sum8[13],carry8[13],sum9[12],carry9[13]);
    full_adder f8_3(k[12],sum9[12],carry9[12],sum10[11],carry10[12]);
    full_adder f8_4(l[11],sum10[11],carry10[11],sum11[10],carry11[11]);
    full_adder f8_5(m[10],sum11[10],carry11[10],sum12[9],carry12[10]);
    full_adder f8_6(n[9],sum12[9],carry12[9],sum13[8],carry13[9]);
    full_adder f8_7(o[8],sum13[8],carry13[8],sum14[7],carry14[8]);
    full_adder f8_8(p[7],sum14[7],carry14[7],sum15[6],carry15[7]);
    full_adder f8_9(sum15[6],carry15[6],carry16[5],out1[22],carry16[6]);

    full_adder f7_1(i[15],j[14],carry8[14],sum9[13],carry9[14]);
    full_adder f7_2(k[13],sum9[13],carry9[13],sum10[12],carry10[13]);
    full_adder f7_3(l[12],sum10[12],carry10[12],sum11[11],carry11[12]);
    full_adder f7_4(m[11],sum11[11],carry11[11],sum12[10],carry12[11]);
    full_adder f7_5(n[10],sum12[10],carry12[10],sum13[9],carry13[10]);
    full_adder f7_6(o[9],sum13[9],carry13[9],sum14[8],carry14[9]);
    full_adder f7_7(p[8],sum14[8],carry14[8],sum15[7],carry15[8]);
    full_adder f7_8(sum15[7],carry15[7],carry16[6],out1[23],carry16[7]);

    full_adder f6_1(j[15],k[14],carry9[14],sum10[13],carry10[14]);
    full_adder f6_2(l[13],sum10[13],carry10[13],sum11[12],carry11[13]);
    full_adder f6_3(m[12],sum11[12],carry11[12],sum12[11],carry12[12]);
    full_adder f6_4(n[11],sum12[11],carry12[11],sum13[10],carry13[11]);
    full_adder f6_5(o[10],sum13[10],carry13[10],sum14[9],carry14[10]);
    full_adder f6_6(p[9],sum14[9],carry14[9],sum15[8],carry15[9]);
    full_adder f6_7(sum15[8],carry15[8],carry16[7],out1[24],carry16[8]);

    full_adder f5_1(k[15],l[14],carry10[14],sum11[13],carry11[14]);
    full_adder f5_2(m[13],sum11[13],carry11[13],sum12[12],carry12[13]);
    full_adder f5_3(n[12],sum12[12],carry12[12],sum13[11],carry13[12]);
    full_adder f5_4(o[11],sum13[11],carry13[11],sum14[10],carry14[11]);
    full_adder f5_5(p[10],sum14[10],carry14[10],sum15[9],carry15[10]);
    full_adder f5_6(sum15[9],carry15[9],carry16[8],out1[25],carry16[9]);

    full_adder f4_1(l[15],m[14],carry11[14],sum12[13],carry12[14]);
    full_adder f4_2(n[13],sum12[13],carry12[13],sum13[12],carry13[13]);
    full_adder f4_3(o[12],sum13[12],carry13[12],sum14[11],carry14[12]);
    full_adder f4_4(p[11],sum14[11],carry14[11],sum15[10],carry15[11]);
    full_adder f4_5(sum15[10],carry15[10],carry16[9],out1[26],carry16[10]);

    full_adder f3_1(m[15],n[14],carry12[14],sum13[13],carry13[14]);
    full_adder f3_2(o[13],sum13[13],carry13[13],sum14[12],carry14[13]);
    full_adder f3_3(p[12],sum14[12],carry14[12],sum15[11],carry15[12]);
    full_adder f3_4(sum15[11],carry15[11],carry16[10],out1[27],carry16[11]);

    full_adder f2_1(n[15],o[14],carry13[14],sum14[13],carry14[14]);
    full_adder f2_2(p[13],sum14[13],carry14[13],sum15[12],carry15[13]);
    full_adder f2_3(sum15[12],carry15[12],carry16[11],out1[28],carry16[12]);

    full_adder f1_1(o[15],p[14],carry14[14],sum15[13],carry15[14]);
    full_adder f1_2(sum15[13],carry15[13],carry16[12],out1[29],carry16[13]);

    full_adder f0_1(p[15],carry15[14],carry16[13],out1[30],out1[31]);

endmodule