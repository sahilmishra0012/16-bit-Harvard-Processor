module shift(a,k);

input  [31:0] a;
//input  [15:0] b;
output [31:0] k;


assign k[0]=0;
assign k[1]=a[0];
assign k[2]=a[1];
assign k[3]=a[2];
assign k[4]=a[3];
assign k[5]=a[4];
assign k[6]=a[5];
assign k[7]=a[6];
assign k[8]=a[7];
assign k[9]=a[8];
assign k[10]=a[9];
assign k[11]=a[10];
assign k[12]=a[11];
assign k[13]=a[12];
assign k[14]=a[13];
assign k[15]=a[14];
assign k[16]=a[15];
assign k[17]=a[16];
assign k[18]=a[17];
assign k[19]=a[18];
assign k[20]=a[19];
assign k[21]=a[20];
assign k[22]=a[21];
assign k[23]=a[22];
assign k[24]=a[23];
assign k[25]=a[24];
assign k[26]=a[25];
assign k[27]=a[26];
assign k[28]=a[27];
assign k[29]=a[28];
assign k[30]=a[29];
assign k[31]=a[30];



/*assign k[32]=a[32];
assign k[33]=a[33];
assign k[34]=a[34];
assign k[35]=a[35];
assign k[36]=a[36];
assign k[37]=a[37];
assign k[38]=a[38];
assign k[39]=a[39];
assign k[40]=a[40];
assign k[41]=a[41];
assign k[42]=a[42];
assign k[43]=a[43];
assign k[44]=a[44];
assign k[45]=a[45];
assign k[46]=a[46];
assign k[47]=a[47];
assign k[48]=a[48];
assign k[49]=a[49];
assign k[50]=a[50];
assign k[51]=a[51];
assign k[52]=a[52];
assign k[53]=a[53];
assign k[54]=a[54];
assign k[55]=a[55];
assign k[56]=a[56];
assign k[57]=a[57];
assign k[58]=a[58];
assign k[59]=a[59];
assign k[60]=a[60];
assign k[61]=a[61];
assign k[62]=a[62];
assign k[63]=a[63];
assign k[64]=a[64];
assign k[65]=a[65];
*/


endmodule
