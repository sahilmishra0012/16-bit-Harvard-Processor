module memory(address,out,read);
input [4:0] address;
output reg [15:0] out;
input read;
reg [15:0] memory [255:0];					
initial
begin
	memory[0]=16'd0;
	memory[1]=16'd1;
	memory[2]=16'd2;
	memory[3]=16'd3;
	memory[4]=16'd4;
	memory[5]=16'd5;
	memory[6]=16'd6;
	memory[7]=16'd7;
	memory[8]=16'd8;
	memory[9]=16'd9;
	memory[10]=16'd10;
	memory[11]=16'd11;
	memory[12]=16'd12;
	memory[13]=16'd13;
	memory[14]=16'd14;
	memory[15]=16'd15;
	memory[16]=16'd16;
	memory[17]=16'd17;
	memory[18]=16'd18;
	memory[19]=16'd19;
	memory[20]=16'd20;
	memory[21]=16'd21;
	memory[22]=16'd22;
	memory[23]=16'd23;
	memory[24]=16'd24;
	memory[25]=16'd25;
	memory[26]=16'd26;
	memory[27]=16'd27;
	memory[28]=16'd28;
	memory[29]=16'd29;
	memory[30]=16'd30;
	memory[31]=16'd31;
	memory[32]=16'd32;
	memory[33]=16'd33;
	memory[34]=16'd34;
	memory[35]=16'd35;
	memory[36]=16'd36;
	memory[37]=16'd37;
	memory[38]=16'd38;
	memory[39]=16'd39;
	memory[40]=16'd40;
	memory[41]=16'd41;
	memory[42]=16'd42;
	memory[43]=16'd43;
	memory[44]=16'd44;
	memory[45]=16'd45;
	memory[46]=16'd46;
	memory[47]=16'd47;
	memory[48]=16'd48;
	memory[49]=16'd49;
	memory[50]=16'd50;
	memory[51]=16'd51;
	memory[52]=16'd52;
	memory[53]=16'd53;
	memory[54]=16'd54;
	memory[55]=16'd55;
	memory[56]=16'd56;
	memory[57]=16'd57;
	memory[58]=16'd58;
	memory[59]=16'd59;
	memory[60]=16'd60;
	memory[61]=16'd61;
	memory[62]=16'd62;
	memory[63]=16'd63;
	memory[64]=16'd64;
	memory[65]=16'd65;
	memory[66]=16'd66;
	memory[67]=16'd67;
	memory[68]=16'd68;
	memory[69]=16'd69;
	memory[70]=16'd70;
	memory[71]=16'd71;
	memory[72]=16'd72;
	memory[73]=16'd73;
	memory[74]=16'd74;
	memory[75]=16'd75;
	memory[76]=16'd76;
	memory[77]=16'd77;
	memory[78]=16'd78;
	memory[79]=16'd79;
	memory[80]=16'd80;
	memory[81]=16'd81;
	memory[82]=16'd82;
	memory[83]=16'd83;
	memory[84]=16'd84;
	memory[85]=16'd85;
	memory[86]=16'd86;
	memory[87]=16'd87;
	memory[88]=16'd88;
	memory[89]=16'd89;
	memory[90]=16'd90;
	memory[91]=16'd91;
	memory[92]=16'd92;
	memory[93]=16'd93;
	memory[94]=16'd94;
	memory[95]=16'd95;
	memory[96]=16'd96;
	memory[97]=16'd97;
	memory[98]=16'd98;
	memory[99]=16'd99;
	memory[100]=16'd100;
	memory[101]=16'd101;
	memory[102]=16'd102;
	memory[103]=16'd103;
	memory[104]=16'd104;
	memory[105]=16'd105;
	memory[106]=16'd106;
	memory[107]=16'd107;
	memory[108]=16'd108;
	memory[109]=16'd109;
	memory[110]=16'd110;
	memory[111]=16'd111;
	memory[112]=16'd112;
	memory[113]=16'd113;
	memory[114]=16'd114;
	memory[115]=16'd115;
	memory[116]=16'd116;
	memory[117]=16'd117;
	memory[118]=16'd118;
	memory[119]=16'd119;
	memory[120]=16'd120;
	memory[121]=16'd121;
	memory[122]=16'd122;
	memory[123]=16'd123;
	memory[124]=16'd124;
	memory[125]=16'd125;
	memory[126]=16'd126;
	memory[127]=16'd127;
	memory[128]=16'd128;
	memory[129]=16'd129;
	memory[130]=16'd130;
	memory[131]=16'd131;
	memory[132]=16'd132;
	memory[133]=16'd133;
	memory[134]=16'd134;
	memory[135]=16'd135;
	memory[136]=16'd136;
	memory[137]=16'd137;
	memory[138]=16'd138;
	memory[139]=16'd139;
	memory[140]=16'd140;
	memory[141]=16'd141;
	memory[142]=16'd142;
	memory[143]=16'd143;
	memory[144]=16'd144;
	memory[145]=16'd145;
	memory[146]=16'd146;
	memory[147]=16'd147;
	memory[148]=16'd148;
	memory[149]=16'd149;
	memory[150]=16'd150;
	memory[151]=16'd151;
	memory[152]=16'd152;
	memory[153]=16'd153;
	memory[154]=16'd154;
	memory[155]=16'd155;
	memory[156]=16'd156;
	memory[157]=16'd157;
	memory[158]=16'd158;
	memory[159]=16'd159;
	memory[160]=16'd160;
	memory[161]=16'd161;
	memory[162]=16'd162;
	memory[163]=16'd163;
	memory[164]=16'd164;
	memory[165]=16'd165;
	memory[166]=16'd166;
	memory[167]=16'd167;
	memory[168]=16'd168;
	memory[169]=16'd169;
	memory[170]=16'd170;
	memory[171]=16'd171;
	memory[172]=16'd172;
	memory[173]=16'd173;
	memory[174]=16'd174;
	memory[175]=16'd175;
	memory[176]=16'd176;
	memory[177]=16'd177;
	memory[178]=16'd178;
	memory[179]=16'd179;
	memory[180]=16'd180;
	memory[181]=16'd181;
	memory[182]=16'd182;
	memory[183]=16'd183;
	memory[184]=16'd184;
	memory[185]=16'd185;
	memory[186]=16'd186;
	memory[187]=16'd187;
	memory[188]=16'd188;
	memory[189]=16'd189;
	memory[190]=16'd190;
	memory[191]=16'd191;
	memory[192]=16'd192;
	memory[193]=16'd193;
	memory[194]=16'd194;
	memory[195]=16'd195;
	memory[196]=16'd196;
	memory[197]=16'd197;
	memory[198]=16'd198;
	memory[199]=16'd199;
	memory[200]=16'd200;
	memory[201]=16'd201;
	memory[202]=16'd202;
	memory[203]=16'd203;
	memory[204]=16'd204;
	memory[205]=16'd205;
	memory[206]=16'd206;
	memory[207]=16'd207;
	memory[208]=16'd208;
	memory[209]=16'd209;
	memory[210]=16'd210;
	memory[211]=16'd211;
	memory[212]=16'd212;
	memory[213]=16'd213;
	memory[214]=16'd214;
	memory[215]=16'd215;
	memory[216]=16'd216;
	memory[217]=16'd217;
	memory[218]=16'd218;
	memory[219]=16'd219;
	memory[220]=16'd220;
	memory[221]=16'd221;
	memory[222]=16'd222;
	memory[223]=16'd223;
	memory[224]=16'd224;
	memory[225]=16'd225;
	memory[226]=16'd226;
	memory[227]=16'd227;
	memory[228]=16'd228;
	memory[229]=16'd229;
	memory[230]=16'd230;
	memory[231]=16'd231;
	memory[232]=16'd232;
	memory[233]=16'd233;
	memory[234]=16'd234;
	memory[235]=16'd235;
	memory[236]=16'd236;
	memory[237]=16'd237;
	memory[238]=16'd238;
	memory[239]=16'd239;
	memory[240]=16'd240;
	memory[241]=16'd241;
	memory[242]=16'd242;
	memory[243]=16'd243;
	memory[244]=16'd244;
	memory[245]=16'd245;
	memory[246]=16'd246;
	memory[247]=16'd247;
	memory[248]=16'd248;
	memory[249]=16'd249;
	memory[250]=16'd250;
	memory[251]=16'd251;
	memory[252]=16'd252;
	memory[253]=16'd253;
	memory[254]=16'd254;
	memory[255]=16'd255;
end


always @(*)

begin

	if(read)
	begin
	out=memory[address];
	end

	else
	begin	
	memory[address]=out;
	out=memory[address];  		
	end

end


endmodule