module and_gate(input [15:0] A,input [15:0] B, output [15:0] OR);
    assign OR = A&B;
endmodule