module left(input [15:0] A, output [15:0] shifted);
    assign shifted = A * 2;
endmodule