module memory(address,out,read);
input [4:0] address;
output reg [15:0] out;
input read;
reg [15:0] memory [255:0];					
initial
begin
	memory[0]=16'b0;
	memory[1]=16'b0;
	memory[2]=16'b0;
	memory[3]=16'b0;
	memory[4]=16'b0;
	memory[5]=16'b0;
	memory[6]=16'b0;
	memory[7]=16'b0;
	memory[8]=16'b0;
	memory[9]=16'b0;
	memory[10]=16'b0;
	memory[11]=16'b0;
	memory[12]=16'b0;
	memory[13]=16'b0;
	memory[14]=16'b0;
	memory[15]=16'b0;
	memory[16]=16'b0;
	memory[17]=16'b0;
	memory[18]=16'b0;
	memory[19]=16'b0;
	memory[20]=16'b0;
	memory[21]=16'b0;
	memory[22]=16'b0;
	memory[23]=16'b0;
	memory[24]=16'b0;
	memory[25]=16'b0;
	memory[26]=16'b0;
	memory[27]=16'b0;
	memory[28]=16'b0;
	memory[29]=16'b0;
	memory[30]=16'b0;
	memory[31]=16'b0;
	memory[32]=16'b0;
	memory[33]=16'b0;
	memory[34]=16'b0;
	memory[35]=16'b0;
	memory[36]=16'b0;
	memory[37]=16'b0;
	memory[38]=16'b0;
	memory[39]=16'b0;
	memory[40]=16'b0;
	memory[41]=16'b0;
	memory[42]=16'b0;
	memory[43]=16'b0;
	memory[44]=16'b0;
	memory[45]=16'b0;
	memory[46]=16'b0;
	memory[47]=16'b0;
	memory[48]=16'b0;
	memory[49]=16'b0;
	memory[50]=16'b0;
	memory[51]=16'b0;
	memory[52]=16'b0;
	memory[53]=16'b0;
	memory[54]=16'b0;
	memory[55]=16'b0;
	memory[56]=16'b0;
	memory[57]=16'b0;
	memory[58]=16'b0;
	memory[59]=16'b0;
	memory[60]=16'b0;
	memory[61]=16'b0;
	memory[62]=16'b0;
	memory[63]=16'b0;
	memory[64]=16'b0;
	memory[65]=16'b0;
	memory[66]=16'b0;
	memory[67]=16'b0;
	memory[68]=16'b0;
	memory[69]=16'b0;
	memory[70]=16'b0;
	memory[71]=16'b0;
	memory[72]=16'b0;
	memory[73]=16'b0;
	memory[74]=16'b0;
	memory[75]=16'b0;
	memory[76]=16'b0;
	memory[77]=16'b0;
	memory[78]=16'b0;
	memory[79]=16'b0;
	memory[80]=16'b0;
	memory[81]=16'b0;
	memory[82]=16'b0;
	memory[83]=16'b0;
	memory[84]=16'b0;
	memory[85]=16'b0;
	memory[86]=16'b0;
	memory[87]=16'b0;
	memory[88]=16'b0;
	memory[89]=16'b0;
	memory[90]=16'b0;
	memory[91]=16'b0;
	memory[92]=16'b0;
	memory[93]=16'b0;
	memory[94]=16'b0;
	memory[95]=16'b0;
	memory[96]=16'b0;
	memory[97]=16'b0;
	memory[98]=16'b0;
	memory[99]=16'b0;
	memory[100]=16'b0;
	memory[101]=16'b0;
	memory[102]=16'b0;
	memory[103]=16'b0;
	memory[104]=16'b0;
	memory[105]=16'b0;
	memory[106]=16'b0;
	memory[107]=16'b0;
	memory[108]=16'b0;
	memory[109]=16'b0;
	memory[110]=16'b0;
	memory[111]=16'b0;
	memory[112]=16'b0;
	memory[113]=16'b0;
	memory[114]=16'b0;
	memory[115]=16'b0;
	memory[116]=16'b0;
	memory[117]=16'b0;
	memory[118]=16'b0;
	memory[119]=16'b0;
	memory[120]=16'b0;
	memory[121]=16'b0;
	memory[122]=16'b0;
	memory[123]=16'b0;
	memory[124]=16'b0;
	memory[125]=16'b0;
	memory[126]=16'b0;
	memory[127]=16'b0;
	memory[128]=16'b0;
	memory[129]=16'b0;
	memory[130]=16'b0;
	memory[131]=16'b0;
	memory[132]=16'b0;
	memory[133]=16'b0;
	memory[134]=16'b0;
	memory[135]=16'b0;
	memory[136]=16'b0;
	memory[137]=16'b0;
	memory[138]=16'b0;
	memory[139]=16'b0;
	memory[140]=16'b0;
	memory[141]=16'b0;
	memory[142]=16'b0;
	memory[143]=16'b0;
	memory[144]=16'b0;
	memory[145]=16'b0;
	memory[146]=16'b0;
	memory[147]=16'b0;
	memory[148]=16'b0;
	memory[149]=16'b0;
	memory[150]=16'b0;
	memory[151]=16'b0;
	memory[152]=16'b0;
	memory[153]=16'b0;
	memory[154]=16'b0;
	memory[155]=16'b0;
	memory[156]=16'b0;
	memory[157]=16'b0;
	memory[158]=16'b0;
	memory[159]=16'b0;
	memory[160]=16'b0;
	memory[161]=16'b0;
	memory[162]=16'b0;
	memory[163]=16'b0;
	memory[164]=16'b0;
	memory[165]=16'b0;
	memory[166]=16'b0;
	memory[167]=16'b0;
	memory[168]=16'b0;
	memory[169]=16'b0;
	memory[170]=16'b0;
	memory[171]=16'b0;
	memory[172]=16'b0;
	memory[173]=16'b0;
	memory[174]=16'b0;
	memory[175]=16'b0;
	memory[176]=16'b0;
	memory[177]=16'b0;
	memory[178]=16'b0;
	memory[179]=16'b0;
	memory[180]=16'b0;
	memory[181]=16'b0;
	memory[182]=16'b0;
	memory[183]=16'b0;
	memory[184]=16'b0;
	memory[185]=16'b0;
	memory[186]=16'b0;
	memory[187]=16'b0;
	memory[188]=16'b0;
	memory[189]=16'b0;
	memory[190]=16'b0;
	memory[191]=16'b0;
	memory[192]=16'b0;
	memory[193]=16'b0;
	memory[194]=16'b0;
	memory[195]=16'b0;
	memory[196]=16'b0;
	memory[197]=16'b0;
	memory[198]=16'b0;
	memory[199]=16'b0;
	memory[200]=16'b0;
	memory[201]=16'b0;
	memory[202]=16'b0;
	memory[203]=16'b0;
	memory[204]=16'b0;
	memory[205]=16'b0;
	memory[206]=16'b0;
	memory[207]=16'b0;
	memory[208]=16'b0;
	memory[209]=16'b0;
	memory[210]=16'b0;
	memory[211]=16'b0;
	memory[212]=16'b0;
	memory[213]=16'b0;
	memory[214]=16'b0;
	memory[215]=16'b0;
	memory[216]=16'b0;
	memory[217]=16'b0;
	memory[218]=16'b0;
	memory[219]=16'b0;
	memory[220]=16'b0;
	memory[221]=16'b0;
	memory[222]=16'b0;
	memory[223]=16'b0;
	memory[224]=16'b0;
	memory[225]=16'b0;
	memory[226]=16'b0;
	memory[227]=16'b0;
	memory[228]=16'b0;
	memory[229]=16'b0;
	memory[230]=16'b0;
	memory[231]=16'b0;
	memory[232]=16'b0;
	memory[233]=16'b0;
	memory[234]=16'b0;
	memory[235]=16'b0;
	memory[236]=16'b0;
	memory[237]=16'b0;
	memory[238]=16'b0;
	memory[239]=16'b0;
	memory[240]=16'b0;
	memory[241]=16'b0;
	memory[242]=16'b0;
	memory[243]=16'b0;
	memory[244]=16'b0;
	memory[245]=16'b0;
	memory[246]=16'b0;
	memory[247]=16'b0;
	memory[248]=16'b0;
	memory[249]=16'b0;
	memory[250]=16'b0;
	memory[251]=16'b0;
	memory[252]=16'b0;
	memory[253]=16'b0;
	memory[254]=16'b0;
	memory[255]=16'b0;
end


always @(*)

begin
	case(read)
	1'b1:
	begin
	out=memory[address];
	end
	1'b0:
	begin	
	memory[address]=out;
	out=memory[address];  		
	end
	endcase
end


endmodule