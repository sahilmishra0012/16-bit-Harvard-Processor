module instruction_set(input );

output [63:0] in [31:0];